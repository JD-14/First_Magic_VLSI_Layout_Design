magic
tech sky130A
timestamp 1634965279
<< nwell >>
rect -332 206 -161 208
rect -332 -15 121 206
rect -163 -17 121 -15
<< nmos >>
rect -251 -183 -236 -141
rect -160 -183 -145 -141
rect 0 -184 15 -142
<< pmos >>
rect -251 14 -236 82
rect -160 14 -145 82
rect 0 14 15 82
<< ndiff >>
rect -300 -154 -251 -141
rect -300 -171 -290 -154
rect -273 -171 -251 -154
rect -300 -183 -251 -171
rect -236 -152 -160 -141
rect -236 -169 -211 -152
rect -194 -169 -160 -152
rect -236 -183 -160 -169
rect -145 -153 -85 -141
rect -145 -170 -133 -153
rect -116 -170 -85 -153
rect -145 -183 -85 -170
rect -55 -142 -38 -141
rect -55 -153 0 -142
rect -55 -170 -28 -153
rect -11 -170 0 -153
rect -55 -183 0 -170
rect -39 -184 0 -183
rect 15 -154 61 -142
rect 15 -171 30 -154
rect 47 -171 61 -154
rect 15 -184 61 -171
<< pdiff >>
rect -306 57 -251 82
rect -306 40 -288 57
rect -271 40 -251 57
rect -306 14 -251 40
rect -236 14 -160 82
rect -145 62 -71 82
rect -145 45 -110 62
rect -93 45 -71 62
rect -145 14 -71 45
rect -43 58 0 82
rect -43 41 -27 58
rect -10 41 0 58
rect -43 14 0 41
rect 15 57 57 82
rect 15 40 27 57
rect 44 40 57 57
rect 15 14 57 40
<< ndiffc >>
rect -290 -171 -273 -154
rect -211 -169 -194 -152
rect -133 -170 -116 -153
rect -28 -170 -11 -153
rect 30 -171 47 -154
<< pdiffc >>
rect -288 40 -271 57
rect -110 45 -93 62
rect -27 41 -10 58
rect 27 40 44 57
<< psubdiff >>
rect -292 -246 -249 -233
rect -292 -263 -280 -246
rect -263 -263 -249 -246
rect -292 -276 -249 -263
rect -195 -245 -152 -232
rect -195 -262 -182 -245
rect -165 -262 -152 -245
rect -195 -275 -152 -262
rect -104 -249 -58 -233
rect -104 -266 -88 -249
rect -70 -266 -58 -249
rect -104 -282 -58 -266
rect 18 -248 61 -231
rect 18 -265 32 -248
rect 49 -265 61 -248
rect 18 -279 61 -265
<< nsubdiff >>
rect -307 147 -264 160
rect -307 130 -294 147
rect -277 130 -264 147
rect -307 117 -264 130
rect -104 145 -54 158
rect -104 128 -88 145
rect -71 128 -54 145
rect -104 113 -54 128
rect 17 144 63 157
rect 17 127 32 144
rect 49 127 63 144
rect 17 114 63 127
<< psubdiffcont >>
rect -280 -263 -263 -246
rect -182 -262 -165 -245
rect -88 -266 -70 -249
rect 32 -265 49 -248
<< nsubdiffcont >>
rect -294 130 -277 147
rect -88 128 -71 145
rect 32 127 49 144
<< poly >>
rect -251 82 -236 101
rect -160 82 -145 100
rect 0 82 15 100
rect -251 -90 -236 14
rect -160 -33 -145 14
rect -189 -41 -145 -33
rect 0 -36 15 14
rect -189 -58 -180 -41
rect -163 -58 -145 -41
rect -189 -67 -145 -58
rect -280 -97 -236 -90
rect -280 -114 -272 -97
rect -255 -114 -236 -97
rect -280 -120 -236 -114
rect -251 -141 -236 -120
rect -160 -141 -145 -67
rect -42 -50 15 -36
rect -42 -67 -31 -50
rect -14 -67 15 -50
rect -42 -84 15 -67
rect 0 -142 15 -84
rect -251 -198 -236 -183
rect -160 -198 -145 -183
rect 0 -200 15 -184
<< polycont >>
rect -180 -58 -163 -41
rect -272 -114 -255 -97
rect -31 -67 -14 -50
<< locali >>
rect -319 147 119 162
rect -319 130 -294 147
rect -277 145 119 147
rect -277 130 -88 145
rect -319 128 -88 130
rect -71 144 119 145
rect -71 128 32 144
rect -319 127 32 128
rect 49 127 119 144
rect -319 113 119 127
rect -300 57 -261 113
rect -150 112 119 113
rect -37 90 -2 112
rect -300 40 -288 57
rect -271 40 -261 57
rect -300 29 -261 40
rect -120 62 -83 71
rect -120 45 -110 62
rect -93 45 -83 62
rect -330 -41 -159 -32
rect -330 -58 -180 -41
rect -163 -58 -159 -41
rect -330 -66 -159 -58
rect -120 -41 -83 45
rect -37 58 -1 90
rect -37 41 -27 58
rect -10 41 -1 58
rect -37 4 -1 41
rect 18 57 54 84
rect 18 40 27 57
rect 44 40 54 57
rect 18 0 54 40
rect -120 -50 -6 -41
rect -120 -67 -31 -50
rect -14 -67 -6 -50
rect -120 -77 -6 -67
rect -330 -97 -245 -89
rect -120 -90 -86 -77
rect -330 -114 -272 -97
rect -255 -114 -245 -97
rect -330 -122 -245 -114
rect -221 -117 -86 -90
rect -298 -154 -264 -142
rect -298 -171 -290 -154
rect -273 -171 -264 -154
rect -298 -225 -264 -171
rect -221 -152 -184 -117
rect -120 -119 -86 -117
rect -221 -169 -211 -152
rect -194 -169 -184 -152
rect -221 -177 -184 -169
rect -143 -153 -105 -143
rect -143 -170 -133 -153
rect -116 -170 -105 -153
rect -143 -225 -105 -170
rect -37 -153 -1 -132
rect -37 -170 -28 -153
rect -11 -170 -1 -153
rect -37 -225 -1 -170
rect 18 -154 53 0
rect 18 -171 30 -154
rect 47 -171 53 -154
rect 18 -194 53 -171
rect -302 -245 120 -225
rect -302 -246 -182 -245
rect -302 -263 -280 -246
rect -263 -262 -182 -246
rect -165 -248 120 -245
rect -165 -249 32 -248
rect -165 -262 -88 -249
rect -263 -263 -88 -262
rect -302 -266 -88 -263
rect -70 -265 32 -249
rect 49 -265 120 -248
rect -70 -266 120 -265
rect -302 -287 120 -266
rect -151 -288 120 -287
<< labels >>
rlabel locali 33 -59 33 -59 1 output
rlabel locali -98 -58 -98 -58 1 n0
rlabel locali -318 -47 -318 -47 1 A
rlabel locali -317 -104 -317 -104 1 B
rlabel locali -25 -255 -25 -255 1 gnd
rlabel locali -22 137 -22 137 1 vdd
rlabel pdiff -202 53 -202 53 1 n1
<< end >>
