magic
tech sky130A
timestamp 1634957434
<< nwell >>
rect -163 -17 121 206
<< nmos >>
rect 0 -184 15 -142
<< pmos >>
rect 0 14 15 82
<< ndiff >>
rect -39 -153 0 -142
rect -39 -170 -28 -153
rect -11 -170 0 -153
rect -39 -184 0 -170
rect 15 -154 61 -142
rect 15 -171 30 -154
rect 47 -171 61 -154
rect 15 -184 61 -171
<< pdiff >>
rect -43 58 0 82
rect -43 41 -27 58
rect -10 41 0 58
rect -43 14 0 41
rect 15 57 57 82
rect 15 40 27 57
rect 44 40 57 57
rect 15 14 57 40
<< ndiffc >>
rect -28 -170 -11 -153
rect 30 -171 47 -154
<< pdiffc >>
rect -27 41 -10 58
rect 27 40 44 57
<< psubdiff >>
rect -104 -249 -58 -233
rect -104 -266 -88 -249
rect -70 -266 -58 -249
rect -104 -282 -58 -266
rect 18 -248 61 -231
rect 18 -265 32 -248
rect 49 -265 61 -248
rect 18 -279 61 -265
<< nsubdiff >>
rect -104 145 -54 158
rect -104 128 -88 145
rect -71 128 -54 145
rect -104 113 -54 128
rect 17 144 63 157
rect 17 127 32 144
rect 49 127 63 144
rect 17 114 63 127
<< psubdiffcont >>
rect -88 -266 -70 -249
rect 32 -265 49 -248
<< nsubdiffcont >>
rect -88 128 -71 145
rect 32 127 49 144
<< poly >>
rect 0 82 15 100
rect 0 -36 15 14
rect -42 -50 15 -36
rect -42 -67 -31 -50
rect -14 -67 15 -50
rect -42 -84 15 -67
rect 0 -142 15 -84
rect 0 -200 15 -184
<< polycont >>
rect -31 -67 -14 -50
<< locali >>
rect -150 145 119 162
rect -150 128 -88 145
rect -71 144 119 145
rect -71 128 32 144
rect -150 127 32 128
rect 49 127 119 144
rect -150 112 119 127
rect -37 90 -2 112
rect -37 58 -1 90
rect -37 41 -27 58
rect -10 41 -1 58
rect -37 4 -1 41
rect 18 57 54 84
rect 18 40 27 57
rect 44 40 54 57
rect 18 0 54 40
rect -54 -50 -6 -41
rect -54 -67 -31 -50
rect -14 -67 -6 -50
rect -54 -77 -6 -67
rect -37 -153 -1 -132
rect -37 -170 -28 -153
rect -11 -170 -1 -153
rect -37 -225 -1 -170
rect 18 -154 53 0
rect 18 -171 30 -154
rect 47 -171 53 -154
rect 18 -194 53 -171
rect -151 -248 120 -225
rect -151 -249 32 -248
rect -151 -266 -88 -249
rect -70 -265 32 -249
rect 49 -265 120 -248
rect -70 -266 120 -265
rect -151 -288 120 -266
<< labels >>
rlabel polycont -23 -58 -23 -58 1 A
rlabel locali 34 -58 34 -58 1 Y
rlabel locali -19 -253 -19 -253 1 gnd
rlabel locali -24 139 -24 139 1 vdd
<< end >>
