magic
tech sky130A
timestamp 1634965423
<< nwell >>
rect -526 206 -161 207
rect -526 -17 121 206
<< nmos >>
rect -392 -185 -377 -143
rect -315 -185 -300 -143
rect 0 -184 15 -142
<< pmos >>
rect -392 14 -377 82
rect -315 14 -300 82
rect 0 14 15 82
<< ndiff >>
rect -443 -154 -392 -143
rect -443 -171 -429 -154
rect -412 -171 -392 -154
rect -443 -185 -392 -171
rect -377 -185 -315 -143
rect -300 -156 -243 -143
rect -300 -173 -277 -156
rect -260 -173 -243 -156
rect -300 -185 -243 -173
rect -39 -153 0 -142
rect -39 -170 -28 -153
rect -11 -170 0 -153
rect -39 -184 0 -170
rect 15 -154 61 -142
rect 15 -171 30 -154
rect 47 -171 61 -154
rect 15 -184 61 -171
<< pdiff >>
rect -450 58 -392 82
rect -450 41 -431 58
rect -414 41 -392 58
rect -450 14 -392 41
rect -377 58 -315 82
rect -377 41 -354 58
rect -337 41 -315 58
rect -377 14 -315 41
rect -300 59 -250 82
rect -300 42 -280 59
rect -263 42 -250 59
rect -300 14 -250 42
rect -43 58 0 82
rect -43 41 -27 58
rect -10 41 0 58
rect -43 14 0 41
rect 15 57 57 82
rect 15 40 27 57
rect 44 40 57 57
rect 15 14 57 40
<< ndiffc >>
rect -429 -171 -412 -154
rect -277 -173 -260 -156
rect -28 -170 -11 -153
rect 30 -171 47 -154
<< pdiffc >>
rect -431 41 -414 58
rect -354 41 -337 58
rect -280 42 -263 59
rect -27 41 -10 58
rect 27 40 44 57
<< psubdiff >>
rect -448 -245 -400 -229
rect -448 -262 -432 -245
rect -415 -262 -400 -245
rect -448 -280 -400 -262
rect -104 -249 -58 -233
rect -104 -266 -88 -249
rect -70 -266 -58 -249
rect -104 -282 -58 -266
rect 18 -248 61 -231
rect 18 -265 32 -248
rect 49 -265 61 -248
rect 18 -279 61 -265
<< nsubdiff >>
rect -449 143 -391 155
rect -449 126 -430 143
rect -413 126 -391 143
rect -449 114 -391 126
rect -300 144 -242 156
rect -300 127 -280 144
rect -263 127 -242 144
rect -300 115 -242 127
rect -104 145 -54 158
rect -104 128 -88 145
rect -71 128 -54 145
rect -104 113 -54 128
rect 17 144 63 157
rect 17 127 32 144
rect 49 127 63 144
rect 17 114 63 127
<< psubdiffcont >>
rect -432 -262 -415 -245
rect -88 -266 -70 -249
rect 32 -265 49 -248
<< nsubdiffcont >>
rect -430 126 -413 143
rect -280 127 -263 144
rect -88 128 -71 145
rect 32 127 49 144
<< poly >>
rect -392 82 -377 96
rect -315 82 -300 97
rect 0 82 15 100
rect -392 -24 -377 14
rect -426 -41 -377 -24
rect -426 -58 -415 -41
rect -398 -58 -377 -41
rect -426 -75 -377 -58
rect -392 -143 -377 -75
rect -315 -77 -300 14
rect 0 -36 15 14
rect -352 -98 -300 -77
rect -42 -50 15 -36
rect -42 -67 -31 -50
rect -14 -67 15 -50
rect -42 -84 15 -67
rect -352 -115 -338 -98
rect -321 -115 -300 -98
rect -352 -128 -300 -115
rect -315 -143 -300 -128
rect 0 -142 15 -84
rect -392 -198 -377 -185
rect -315 -200 -300 -185
rect 0 -200 15 -184
<< polycont >>
rect -415 -58 -398 -41
rect -31 -67 -14 -50
rect -338 -115 -321 -98
<< locali >>
rect -518 145 119 162
rect -518 144 -88 145
rect -518 143 -280 144
rect -518 126 -430 143
rect -413 127 -280 143
rect -263 128 -88 144
rect -71 144 119 145
rect -71 128 32 144
rect -263 127 32 128
rect 49 127 119 144
rect -413 126 119 127
rect -518 112 119 126
rect -518 107 -148 112
rect -442 58 -405 107
rect -442 41 -431 58
rect -414 41 -405 58
rect -442 24 -405 41
rect -363 58 -326 70
rect -363 41 -354 58
rect -337 41 -326 58
rect -363 -27 -326 41
rect -290 59 -253 107
rect -290 42 -280 59
rect -263 42 -253 59
rect -290 26 -253 42
rect -37 90 -2 112
rect -37 58 -1 90
rect -37 41 -27 58
rect -10 41 -1 58
rect -37 4 -1 41
rect 18 57 54 84
rect 18 40 27 57
rect 44 40 54 57
rect 18 0 54 40
rect -498 -41 -390 -31
rect -498 -58 -415 -41
rect -398 -58 -390 -41
rect -498 -69 -390 -58
rect -363 -35 -325 -27
rect -363 -39 -252 -35
rect -363 -41 -52 -39
rect -363 -50 -6 -41
rect -363 -65 -31 -50
rect -286 -67 -31 -65
rect -14 -67 -6 -50
rect -286 -76 -6 -67
rect -499 -98 -312 -89
rect -499 -115 -338 -98
rect -321 -115 -312 -98
rect -499 -124 -312 -115
rect -438 -154 -401 -142
rect -438 -171 -429 -154
rect -412 -171 -401 -154
rect -438 -224 -401 -171
rect -286 -156 -252 -76
rect -54 -77 -6 -76
rect -286 -173 -277 -156
rect -260 -173 -252 -156
rect -286 -183 -252 -173
rect -37 -153 -1 -132
rect -37 -170 -28 -153
rect -11 -170 -1 -153
rect -500 -225 -150 -224
rect -37 -225 -1 -170
rect 18 -154 53 0
rect 18 -171 30 -154
rect 47 -171 53 -154
rect 18 -194 53 -171
rect -500 -245 120 -225
rect -500 -262 -432 -245
rect -415 -248 120 -245
rect -415 -249 32 -248
rect -415 -262 -88 -249
rect -500 -266 -88 -262
rect -70 -265 32 -249
rect 49 -265 120 -248
rect -70 -266 120 -265
rect -500 -287 120 -266
rect -151 -288 120 -287
<< labels >>
rlabel locali -183 -254 -183 -254 1 gnd
rlabel locali -181 134 -181 134 1 vdd
rlabel locali -473 -106 -473 -106 1 A
rlabel locali -475 -50 -475 -50 1 B
rlabel locali -151 -60 -151 -60 1 n0
rlabel locali 34 -61 34 -61 1 output
rlabel ndiff -350 -160 -350 -160 1 n1
<< end >>
